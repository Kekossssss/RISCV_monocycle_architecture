//Author : Kevin GUILLOUX
//Last modified : 11/05/2024
//Comment : Package for the RISCV32i architecture

package RISCV32i_Pack;
	typedef logic [31:0] data_bus;
	typedef logic [2:0] funct3;
	typedef logic [6:0] funct7;
	typedef logic [4:0] adresse_registre;
	typedef logic [6:0] opcode;
endpackage : RISCV32i_Pack
